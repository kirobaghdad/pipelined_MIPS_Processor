library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Execution_Stage is
  port (
    -- INPUTS 
    clk : in std_logic;
    rst : in std_logic;
    user_input: in std_logic_vector(15 downto 0);
    R1 : in STD_LOGIC_VECTOR (15 downto 0);
    R2 : in STD_LOGIC_VECTOR (15 downto 0);
    updated_PC : in STD_LOGIC_VECTOR (15 downto 0);
    IMMD : in STD_LOGIC_VECTOR (15 downto 0);
    Rdst : in STD_LOGIC_VECTOR (2 downto 0);

    
    -- Control Signals
    mem_read : in std_logic;
    mem_write : in std_logic;
    reg_write : in std_logic;
    alu_control : in STD_LOGIC_VECTOR (2 downto 0);
    in_control : in STD_LOGIC;
    IMMD_Control : in STD_LOGIC;

    branch : in std_logic;
    mem_to_reg : in std_logic;
    stack : in std_logic;
    call : in std_logic;
    pop : in std_logic;
    ldm: in std_logic;
    ret: in std_logic;
    rti: in std_logic;
    store : in std_logic;
    int : in std_logic;
    zero : in std_logic;
    enable : in std_logic;


    -- Outputs 
    e_reg_write : out std_logic;
    e_Rdst : out std_logic_vector(2 downto 0);
    e_updated_PC : out std_logic_vector(15 downto 0);
    e_result : out std_logic_vector(15 downto 0);
    e_mem_read : out std_logic;
    e_mem_write : out std_logic;

    e_mem_to_reg : out std_logic;
    e_stack : out std_logic;
    e_call : out std_logic;
    e_pop : out std_logic;
    e_ldm: out std_logic;
    e_ret: out std_logic;
    e_rti: out std_logic;
    e_store : out std_logic;
    e_int : out std_logic;
    e_enable : out std_logic
    -- e_IMMD_Control : out STD_LOGIC;
    -- e_zero : out std_logic;
    -- branch : in std_logic;
    
  ) ;
end Execution_Stage;


architecture behavioral of Execution_Stage is
  signal OP1 : std_logic_vector(15 downto 0);
  signal temp_result : std_logic_vector(15 downto 0);
begin
    uut1: entity work.alu PORT MAP(alu_control => alu_control, OP1 => OP1, OP2 => R2, old_CCR => "000", result => temp_result);

    uut2: entity work.Ex_MEM_Reg PORT MAP(clk => clk, rst => rst, reg_write => reg_write, Rdst => Rdst, updated_PC => updated_PC, mem_read => mem_read, mem_write => mem_write, mem_to_reg => mem_to_reg, stack => stack, call => call, pop => pop, ldm => ldm, ret => ret, rti => rti, store => store, int => int, enable => enable, result => temp_result, reg_write_r => e_reg_write, Rdst_r => e_Rdst, updated_PC_r => e_updated_PC, result_r => e_result, mem_read_r => e_mem_read, mem_write_r => e_mem_write, mem_to_reg_r => e_mem_to_reg, stack_r => e_stack, call_r=> e_call, pop_r => e_pop, ldm_r => e_ldm, ret_r => e_ret, rti_r => e_rti, store_r => e_store, int_r => e_int, enable_r => e_enable);

    uut3: entity work.R1_Selector PORT MAP(IMMD_Control => IMMD_Control, in_control => in_control, IMMD => IMMD, user_input => user_input, R1 => R1, OP1 => OP1);
    
    
end architecture behavioral;